`timescale 1ns / 1ps
/////////////////////////////////////////////////////////////////
// Module Name: xup_and2
/////////////////////////////////////////////////////////////////
module xup_and2 #(parameter DELAY=3)(
    input a,
    input b,
    output y
    );

    and #DELAY (y, a, b);

endmodule
